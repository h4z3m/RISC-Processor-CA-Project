-- LIBRARY IEEE
-- LIBRARY work;
-- USE IEEE.std_logic_1164.ALL;
-- USE IEEE.numeric_std.ALL;
-- ENTITY byte_addressable_memory IS
--     PORT (
--         clk : IN STD_LOGIC;
--         rdwr : IN STD_LOGIC;
--         addr : IN unsigned(11 DOWNTO 0);
--         size : IN unsigned(1 DOWNTO 0);
--         idata : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
--         odata : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
--         ivalid : OUT STD_LOGIC
--     );
-- END ENTITY byte_addressable_memory;

-- ARCHITECTURE rtl OF byte_addressable_memory IS
--     TYPE mem_type IS ARRAY (4095 DOWNTO 0) OF STD_LOGIC_VECTOR(31 DOWNTO 0);
--     SIGNAL mem : mem_type := (OTHERS => (OTHERS => '0'));
-- BEGIN
--     PROCESS (clk)
--     BEGIN
--         IF rising_edge(clk) THEN
--             IF rdwr = '1' THEN
--                 CASE size IS
--                     WHEN "00" =>
--                         mem(to_integer(unsigned(addr))) <= idata(7 DOWNTO 0) & mem(to_integer(unsigned(addr)))(31 DOWNTO 8);
--                         mem(to_integer(unsigned(addr)) + 1) <= idata(15 DOWNTO 8) & mem(to_integer(unsigned(addr)) + 1)(31 DOWNTO 16);
--                         mem(to_integer(unsigned(addr)) + 2) <= idata(23 DOWNTO 16) & mem(to_integer(unsigned(addr)) + 2)(31 DOWNTO 24);
--                         mem(to_integer(unsigned(addr)) + 3) <= idata(31 DOWNTO 24) & mem(to_integer(unsigned(addr)) + 3)(31 DOWNTO 24);
--                     WHEN "01" =>
--                         mem(to_integer(unsigned(addr))) <= idata(15 DOWNTO 0) & mem(to_integer(unsigned(addr)))(31 DOWNTO 16);
--                         mem(to_integer(unsigned(addr)) + 1) <= idata(31 DOWNTO 16) & mem(to_integer(unsigned(addr)) + 1)(31 DOWNTO 16);
--                     WHEN OTHERS =>
--                         NULL;
--                 END CASE;
--                 -- Wait for write to complete
--                 FOR i IN 1 TO 8 LOOP
--                     IF i = 8 THEN
--                         -- Writing complete
--                         ivalid <= '0';
--                     ELSE
--                         -- Writing still in progress
--                         ivalid <= '1';
--                     END IF;
--                     WAIT UNTIL rising_edge(clk);
--                 END LOOP;
--             ELSE
--                 CASE size IS
--                     WHEN "00" =>
--                         odata <= mem(to_integer(unsigned(addr)));
--                     WHEN "01" =>
--                         odata <= mem(to_integer(unsigned(addr)));
--                         odata(15 DOWNTO 0) <= (OTHERS => 'Z');
--                     WHEN OTHERS =>
--                         NULL;
--                 END CASE;
--             END IF;
--         END IF;
--     END PROCESS;
-- END ARCHITECTURE rtl