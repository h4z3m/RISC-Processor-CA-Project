LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;
LIBRARY work;
LIBRARY work;
ENTITY ALU IS
    PORT (
        Opcode : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
        Operand_1 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        Operand_2 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        Output : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
        CARRY : OUT STD_LOGIC;
        ZERO : OUT STD_LOGIC;
        NEGATIVE : OUT STD_LOGIC
    );
END ENTITY ALU;